module ram(i_clk, i_addr, i_data, i_we, o_data);
parameter DATA_WIDTH = 32;
parameter ADDR_WIDTH = 5; //32 4-byte words 

input                     i_clk, i_we;
input   [ADDR_WIDTH-1:0]  i_addr;
input   [DATA_WIDTH-1:0]  i_data;
output  [DATA_WIDTH-1:0]  o_data;

reg	[DATA_WIDTH-1:0]	m_ram[0:(2**ADDR_WIDTH)-1];

initial begin
$readmemh("ram_init.dat", m_ram);
end


always @(posedge i_clk) begin
	if(i_we) begin
		m_ram[i_addr] = i_data;
		$writememh("Debug/ram_result.dat", m_ram);
	end
end
  
assign o_data = m_ram[i_addr];

endmodule
